module MAC(input [71:0] image, 
           input [35:0] weight, 
           input [4:0] exp_bias, 
           output reg [15:0] out);

    


    always @ (image or weight or exp_bias) begin
        
    end
        


endmodule